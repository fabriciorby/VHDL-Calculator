LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;
USE IEEE.NUMERIC_STD.all;


ENTITY CALCULADORA IS
	PORT ( 

		------------------------	Clock Input	 	------------------------
		CLOCK_24	: 	IN	STD_LOGIC_VECTOR (1 DOWNTO 0);	--	24 MHz
		CLOCK_27	:	IN	STD_LOGIC_VECTOR (1 DOWNTO 0);	--	27 MHz
		CLOCK_50	: 	IN	STD_LOGIC;						--	50 MHz
		
		------------------------	Push Button		------------------------
		KEY 	:		IN	STD_LOGIC_VECTOR (3 DOWNTO 0);		--	PUSHBUTTON[3:0]

		------------------------	DPDT Switch		------------------------
		SW 		:		IN STD_LOGIC_VECTOR (9 DOWNTO 0);			--	TOGGLE SWITCH[9:0]
		
		------------------------	7-SEG Display	------------------------
		HEX0 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	SEVEN SEGMENT DIGIT 0
		HEX1 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	SEVEN SEGMENT DIGIT 1
		HEX2 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	SEVEN SEGMENT DIGIT 2
		HEX3 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	Seven Segment Digit 3
		
		----------------------------	LED		----------------------------
		LEDG 	:		OUT	STD_LOGIC_VECTOR (7 DOWNTO 0);		--	LED GREEN[7:0]
		LEDR 	:		OUT	STD_LOGIC_VECTOR (9 DOWNTO 0);		--	LED Red[9:0]
					
		------------------------	PS2		--------------------------------
		PS2_DAT :		INOUT	STD_LOGIC;	--	PS2 Data
		PS2_CLK	:		INOUT	STD_LOGIC	--	PS2 Clock
	);

END CALCULADORA;

ARCHITECTURE funcionamento OF CALCULADORA IS
			
	-- IMPORTANDO COMPONENTES --

	-- CONTROLADOR DE BRILHO DO DISPLAY
	COMPONENT PWM 
		PORT ( 
			CLOCK	: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			ENABLE	: IN STD_LOGIC;
			DUTY	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			CIN		: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			COUTP	: BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0)
		);
	END COMPONENT;

	-- CONVERSOR DE SCANCODE PARA VALOR DE ENTRADA
	COMPONENT conv_calc
		PORT (
			SCAN	:		IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			ENTRADA	:		OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
		);
	END COMPONENT;

	-- CONVERSOR PARA 7SEG
	COMPONENT conv_7seg
		PORT (
			DIGIT	:		IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			SEG		:		OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		);
	END COMPONENT;

	-- BINARY TO BCD
	COMPONENT binary_to_bcd
    	PORT (
			BINARY 		: IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
           	BCD_UNI 	: OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
           	BCD_TEN 	: OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
           	BCD_HUN 	: OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
           	BCD_THO 	: OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
        );
	END COMPONENT;
	
	-- SOMADOR BINARIO PARALELO (NÃO INTEGRADO)

	-- COMPONENT testaSomador
	-- 	GENERIC (N : INTEGER);
	-- 	PORT( 
	-- 		A, B	: IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
	-- 		S		: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0);
	-- 		COUT	: OUT STD_LOGIC
	-- 	);
	-- END COMPONENT;

	-- BIBLIOTECA PARA CONTROLE DO TECLADO
	COMPONENT kbdex_ctrl
		GENERIC (
			CLKFREQ : INTEGER
		);
		PORT (
			PS2_DATA	:	INOUT STD_LOGIC;
			PS2_CLK		:	INOUT STD_LOGIC;
			CLK			:	IN STD_LOGIC;
			EN			:	IN STD_LOGIC;
			RESETN		:	IN STD_LOGIC;
			LIGHTS		:	IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- LIGHTS(CAPS, NUN, SCROLL)		
			KEY_ON		:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
			KEY_CODE	:	OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
		);
	END COMPONENT;
	
	-- DECLARACAO DE SIGNALS
		
	SIGNAL COUT 	: STD_LOGIC := '0';
	SIGNAL COUTP 	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL DUTY	: 	 STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL ENTRADA 	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL BINARY 	: STD_LOGIC_VECTOR (11 DOWNTO 0);
	SIGNAL DIGITOS 	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL RESETN	: STD_LOGIC;
	SIGNAL RESET	: STD_LOGIC;
	SIGNAL key0 	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL lights	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL key_on	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL key_code	: STD_LOGIC_VECTOR (47 DOWNTO 0);

	-- CONSTANTES DEFINIDAS EM conv_calc.vhd

	CONSTANT SUM : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1010"; -- SOMA
	CONSTANT SUB : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1011"; -- SUBTRAÇÃO
	CONSTANT MUL : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1100"; -- MULTIPLICAÇÃO
	CONSTANT DIV : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1101"; -- DIVISÃO
	CONSTANT ENT : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1110"; -- ENTER
	CONSTANT BKS : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1111";	-- BACKSPACE

	CONSTANT VAZIO : STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');

	BEGIN

	-- PROCESS

	PROCESS(ENTRADA, RESET, KEY_ON(0))

	VARIABLE COUNT  : INTEGER := 0;
	VARIABLE OP		: INTEGER := 0;
	VARIABLE A 		: STD_LOGIC_VECTOR (11 DOWNTO 0) := VAZIO;
	VARIABLE B 		: STD_LOGIC_VECTOR (11 DOWNTO 0) := VAZIO;
	VARIABLE C 		: STD_LOGIC_VECTOR (11 DOWNTO 0) := VAZIO;
	VARIABLE D 		: STD_LOGIC_VECTOR (11 DOWNTO 0) := VAZIO;
	VARIABLE TEMP	: STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');

	BEGIN
		IF (RESET = '0') THEN 
			BINARY <= VAZIO;
			A:=VAZIO;
			B:=VAZIO;
			C:=VAZIO;
			D:=VAZIO;
			OP:= 0;
			COUT <= '0';
		ELSIF (key_on(0)'EVENT AND key_on(0) = '1') THEN
					
			CASE ENTRADA IS

				WHEN SUM =>

					COUNT := 0;
					OP := 1;

					IF (A = VAZIO) THEN 
						A := BINARY;
						C := A;
						B := VAZIO;
					END IF;

				WHEN SUB =>

					COUNT := 0;
					OP := 2;

					IF (A = VAZIO) THEN 
						A := BINARY;
						C := A;
						B := VAZIO;
					END IF;

				WHEN MUL =>

					COUNT := 0;
					OP := 3;

					-- CÓDIGO DE MULTIPLICAÇÃO DELETADO

				WHEN DIV =>

					COUNT := 0;
					OP := 4;

					-- CÓDIGO DE DIVISÃO DELETADO

				WHEN ENT =>

					COUNT := 0;

					IF (B = VAZIO) THEN
						B := BINARY;
					END IF;
					
					CASE OP IS 
							WHEN 1 =>
								D := C + BINARY;
								IF (C(11) = '0') AND (BINARY(11) = '0') THEN 
									IF D(11) = '1' THEN
										COUT <= '1'; -- OVERFLOW
									END IF;
								END IF;
								BINARY <= C + BINARY;
								C := B;
							WHEN 2 =>
								D := C - B;
								IF (C(11) = '1') AND (B(11) = '0') THEN 
									IF D(11) = '0' THEN
										COUT <= '1'; -- UNDERFLOW
									END IF;
								END IF;
								BINARY <= C - B;
								C := C - B;
							WHEN 3 =>
								-- CÓDIGO DE MULTIPLICAÇÃO DELETADO
							WHEN 4 =>
								-- CÓDIGO DE DIVISÃO DELETADO
							WHEN OTHERS =>
					END CASE;
					
					A := VAZIO;
					
				WHEN BKS =>
					-- CÓDIGO DE BACKSPACE NECESSITA DA DIVISÃO POR 10

					-- IF NOT (COUNT = 0) THEN
						-- BINARY <= BINARY/10;
						-- COUNT := COUNT - 1;
					-- END IF;
				WHEN OTHERS =>
					IF NOT (BINARY = VAZIO AND ENTRADA = "0000") THEN
						CASE COUNT IS
							WHEN 0 =>
								BINARY <= VAZIO + ENTRADA;
								COUNT := COUNT + 1;
							WHEN 1 TO 3 =>
								D := BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + ENTRADA;
								IF (D(11) = '1') THEN 
									COUT <= '1'; -- OVERFLOW
								END IF;
								BINARY <= BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + BINARY + ENTRADA;
								COUNT := COUNT + 1;
							WHEN OTHERS =>
						END CASE;
					END IF;
			END CASE;
		END IF;
	END PROCESS;

	DUTY	<= SW(7 DOWNTO 0);
	
	RESETN <= KEY(0);
	
	RESET <= KEY(1);
	
	--PEGA OS CLIQUES DO TECLADO

	kbd_ctrl : kbdex_ctrl GENERIC MAP(24000) PORT MAP(
		PS2_DAT, PS2_CLK, CLOCK_24(0), KEY(1), resetn, lights,
		key_on, key_code(15 DOWNTO 0) => key0
	);

	--TRANSFORMA OS CLIQUES EM COMANDOS

	dig_calc: conv_calc PORT MAP (
		key0(7 DOWNTO 0), ENTRADA
	);

	-- SOMADOR DE DOIS NÚMEROS BINÁRIOS (NÃO INTEGRADO)

	--somador: testaSomador GENERIC MAP(12) PORT MAP (
	--	A, B,
	--	SOMA, COUT
	--);

	--TRANSFORMA OS NUMEROS BINARIOS EM 4 CASAS DECIMAIS

	bin2bcd: binary_to_bcd PORT MAP (
		BINARY, 	
		DIGITOS (3 DOWNTO 0), DIGITOS (7 DOWNTO 4), DIGITOS (11 DOWNTO 8), DIGITOS (15 DOWNTO 12) 
	);

	--CONTROLA O BRILHO DO DISPLAY DE 7 SEGMENTOS

	controlador: PWM PORT MAP (
		CLOCK_50,
		RESET, 
		RESETN, --KEY(0)
		DUTY, 
		DIGITOS,
		COUTP
	);

	--MOSTRA OS NUMEROS NO DISPLAY DE 7 SEGMENTOS COM BRILHO CONTROLADO

	hexseg0: conv_7seg PORT MAP (
		COUTP (3 DOWNTO 0), HEX0
	);
	hexseg1: conv_7seg PORT MAP (
		COUTP (7 DOWNTO 4), HEX1
	);
	hexseg2: conv_7seg PORT MAP (
		COUTP (11 DOWNTO 8), HEX2
	);
	hexseg3: conv_7seg PORT MAP (
		COUTP (15 DOWNTO 12), HEX3
	);
	
	--CHECA OVERFLOW
	
	WITH COUT SELECT
		LEDR <=  "1111111111" WHEN '1',
				   "0000000000" WHEN '0';
	
	--CHECA NEGATIVO
	
	WITH BINARY(11) SELECT
		LEDG <= 	"11111111" WHEN '1',
					"00000000" WHEN '0';

END funcionamento;