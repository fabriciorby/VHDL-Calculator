library verilog;
use verilog.vl_types.all;
entity somadorCompleto_vlg_vec_tst is
end somadorCompleto_vlg_vec_tst;
