library verilog;
use verilog.vl_types.all;
entity atividadeMoore_vlg_vec_tst is
end atividadeMoore_vlg_vec_tst;
