library verilog;
use verilog.vl_types.all;
entity binary4_to_bcd8_vector_vlg_vec_tst is
end binary4_to_bcd8_vector_vlg_vec_tst;
