LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY TestaSomador IS
	GENERIC (N : INTEGER := 8);
	PORT ( 
		A, B	: IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		S		: BUFFER STD_LOGIC_VECTOR (N-1 DOWNTO 0);
		COUT	: OUT STD_LOGIC
	);

END TestaSomador;

ARCHITECTURE funcionamento OF TestaSomador IS

	COMPONENT somadorBinarioParalelo
		GENERIC (N : INTEGER);
		PORT( 
			A, B	: IN  STD_LOGIC_VECTOR (N-1 DOWNTO 0);
			CIN	: IN  STD_LOGIC;
			S		: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0);
			COUT	: OUT STD_LOGIC
		);
	END COMPONENT;
	
	SIGNAL E : STD_LOGIC_VECTOR (N-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL OVERFLOW : STD_LOGIC;
	
	BEGIN
						
	COUT <= (A(N-1) AND B(N-1) AND NOT(S(N-1))) OR (NOT(A(N-1)) AND NOT(B(N-1)) AND S(N-1));
	
	somador: somadorBinarioParalelo GENERIC MAP(N) PORT MAP (
		A, B, '0',
		S, OVERFLOW
	);
		
END funcionamento;