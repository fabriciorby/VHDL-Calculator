library verilog;
use verilog.vl_types.all;
entity somadorBinarioParalelo_vlg_vec_tst is
end somadorBinarioParalelo_vlg_vec_tst;
