library verilog;
use verilog.vl_types.all;
entity paridade_hierarquico_vlg_check_tst is
    port(
        p               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end paridade_hierarquico_vlg_check_tst;
