library verilog;
use verilog.vl_types.all;
entity maquinaMoore_vlg_vec_tst is
end maquinaMoore_vlg_vec_tst;
