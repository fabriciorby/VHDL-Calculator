library verilog;
use verilog.vl_types.all;
entity somadorCompleto_vlg_check_tst is
    port(
        COUT            : in     vl_logic;
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end somadorCompleto_vlg_check_tst;
