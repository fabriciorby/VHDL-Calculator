library verilog;
use verilog.vl_types.all;
entity divisorDeClock_vlg_vec_tst is
end divisorDeClock_vlg_vec_tst;
