library verilog;
use verilog.vl_types.all;
entity divisorDeClock_vlg_check_tst is
    port(
        COUT            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end divisorDeClock_vlg_check_tst;
