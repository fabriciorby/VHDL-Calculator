library verilog;
use verilog.vl_types.all;
entity maquinaMoore2_vlg_vec_tst is
end maquinaMoore2_vlg_vec_tst;
