library verilog;
use verilog.vl_types.all;
entity paridade_hierarquico_vlg_vec_tst is
end paridade_hierarquico_vlg_vec_tst;
