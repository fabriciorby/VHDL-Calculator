library verilog;
use verilog.vl_types.all;
entity atividadeMoore_vlg_check_tst is
    port(
        z               : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end atividadeMoore_vlg_check_tst;
