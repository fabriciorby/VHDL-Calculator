LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.std_logic_unsigned.all;


ENTITY PWM IS
	PORT ( 
		CLOCK		: IN  STD_LOGIC;
		RESET		: IN  STD_LOGIC;
		ENABLE	: IN  STD_LOGIC;
		DUTY		: IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		CIN		: IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		COUTP		: BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0)
	);

END PWM;

ARCHITECTURE funcionamento OF pwm IS
		
	SIGNAL COUNT : STD_LOGIC_VECTOR (7 DOWNTO 0);
	
	BEGIN
	
	PROCESS (RESET, CLOCK, ENABLE)
										
	BEGIN
							
		IF RESET = '0' THEN
		
			COUNT <= "00000000";
			
			COUTP <= (OTHERS => '1');
			
		ELSIF (ENABLE = '0') THEN
						
			COUTP <= CIN;

		ELSIF (CLOCK'EVENT AND CLOCK = '1') THEN				
			
			COUNT <= COUNT + '1';
			
			IF (COUNT <= DUTY) THEN
			
				COUTP <= CIN;
			
			ELSIF (COUNT = "11111111") THEN
			
				COUNT <= "00000000";
			
			ELSE
			
				COUTP <= (OTHERS => '1');
			
			END IF;
			
		END IF;
		
	END PROCESS;
			
END funcionamento;