LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.std_logic_unsigned.all;


ENTITY CALC IS
	PORT ( 

		-- PWM --
		CLOCK	: IN  STD_LOGIC;
		RESET	: IN  STD_LOGIC;
		ENABLE	: IN  STD_LOGIC;
		DUTY	: IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		COUT	: BUFFER STD_LOGIC

		------------------------	Clock Input	 	------------------------
		CLOCK_24	: 	IN	STD_LOGIC_VECTOR (1 DOWNTO 0);	--	24 MHz
		CLOCK_27	:	IN	STD_LOGIC_VECTOR (1 DOWNTO 0);	--	27 MHz
		CLOCK_50	: 	IN	STD_LOGIC;						--	50 MHz
		-- CLOCKTAP	: 	OUT	STD_LOGIC;
		
		------------------------	Push Button		------------------------
		KEY 	:		IN	STD_LOGIC_VECTOR (3 DOWNTO 0);		--	PUSHBUTTON[3:0]

		------------------------	DPDT Switch		------------------------
		SW 		:		IN STD_LOGIC_VECTOR (9 DOWNTO 0);			--	TOGGLE SWITCH[9:0]
		
		------------------------	7-SEG Display	------------------------
		HEX0 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	SEVEN SEGMENT DIGIT 0
		HEX1 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	SEVEN SEGMENT DIGIT 1
		HEX2 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	SEVEN SEGMENT DIGIT 2
		HEX3 	:		OUT	STD_LOGIC_VECTOR (6 DOWNTO 0);		--	Seven Segment Digit 3
		
		----------------------------	LED		----------------------------
		LEDG 	:		OUT	STD_LOGIC_VECTOR (7 DOWNTO 0);		--	LED GREEN[7:0]
		LEDR 	:		OUT	STD_LOGIC_VECTOR (9 DOWNTO 0);		--	LED Red[9:0]
					
		------------------------	PS2		--------------------------------
		PS2_DAT :		INOUT	STD_LOGIC;	--	PS2 Data
		PS2_CLK	:		INOUT	STD_LOGIC	--	PS2 Clock
	);

END CALC;

ARCHITECTURE funcionamento OF CALC IS
			
	-- IMPORTANDO COMPONENTES --

	-- CONTROLADOR DE BRILHO DO DISPLAY
	COMPONENT PWM 
		PORT ( 
			CLOCK	: IN STD_LOGIC;
			RESET	: IN STD_LOGIC;
			ENABLE	: IN STD_LOGIC;
			DUTY	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			COUT	: BUFFER STD_LOGIC
		);
	END COMPONENT;

	-- CONVERSOR DE SCANCODE PARA VALOR DE ENTRADA
	COMPONENT conv_calc
		PORT (
			SCAN	:		IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			ENTRADA	:		OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		);
	END COMPONENT;

	-- CONVERSOR PARA 7SEG
		COMPONENT conv_7seg
		PORT (
			DIGIT	:		IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			SEG		:		OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
		);
	END COMPONENT;

	-- BIBLIOTECA PARA CONTROLE DO TECLADO
	COMPONENT kbdex_ctrl
		GENERIC (
			CLKFREQ : INTEGER
		);
		PORT (
			PS2_DATA	:	INOUT STD_LOGIC;
			PS2_CLK		:	INOUT STD_LOGIC;
			CLK			:	IN STD_LOGIC;
			EN			:	IN STD_LOGIC;
			RESETN		:	IN STD_LOGIC;
			LIGHTS		:	IN STD_LOGIC_VECTOR(2 DOWNTO 0); -- LIGHTS(CAPS, NUN, SCROLL)		
			KEY_ON		:	OUT	STD_LOGIC_VECTOR(2 DOWNTO 0);
			KEY_CODE	:	OUT	STD_LOGIC_VECTOR(47 DOWNTO 0)
		);
	END COMPONENT;

	-- DECLARACAO DE SIGNALS

	SIGNAL ENTRADA 	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL DIGITOS 	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL DBUFFER 	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL A 		: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL B 		: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL CIN		: STD_LOGIC_VECTOR (3 DOWNTO 0);

	-- CONSTANTES DEFINIDAS EM conv_calc.vhd

	CONSTANT SUM : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1010";
	CONSTANT SUB : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1011";
	CONSTANT MUL : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1100";
	CONSTANT DIV : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1101";
	CONSTANT ENT : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1110";
	CONSTANT BKS : STD_LOGIC_VECTOR (3 DOWNTO 0) := "1111";

	CONSTANT VAZIO : STD_LOGIC_VECTOR (3 DOWNTO 0) := "0000000000000000";

	BEGIN

	-- PROCESS

	PROCESS(ENTRADA)

	VARIABLE COUNT : INTEGER;

	BEGIN

		CASE ENTRADA IS
			WHEN SUM =>

				COUNT := 0;

				IF (A = VAZIO) THEN 
					A := DIGITOS;
					DIGITOS := VAZIO;
				ELSIF (B = VAZIO) THEN
					B := DIGITOS;
					DIGITOS := DBUFFER;
					A := VAZIO;
					B := VAZIO;
				END IF;

			WHEN SUB =>
				COUNT := 0;
				A := DIGITOS;
				DIGITOS := VAZIO;
			WHEN MUL =>
				COUNT := 0;
				A := DIGITOS;
				DIGITOS := VAZIO;
			WHEN DIV =>
				COUNT := 0;
				A := DIGITOS;
				DIGITOS := VAZIO;
			WHEN OTHERS =>
				IF NOT (DIGITOS = VAZIO AND ENTRADA = "0000") THEN
					CASE COUNT IS
						WHEN 0 =>
							DIGITOS (3 DOWNTO 0) = ENTRADA;
							COUNT := COUNT + 1
						WHEN 1 =>
							DIGITOS (7 DOWNTO 4) = DIGITOS (3 DOWNTO 0);
							DIGITOS (3 DOWNTO 0) = ENTRADA;
							COUNT := COUNT + 1
						WHEN 2 =>
							DIGITOS (11 DOWNTO 8) = DIGITOS (7 DOWNTO 4);
							DIGITOS (7 DOWNTO 4) = DIGITOS (3 DOWNTO 0);
							DIGITOS (3 DOWNTO 0) = ENTRADA;
							COUNT := COUNT + 1
						WHEN 3 =>
							DIGITOS (15 DOWNTO 12) = DIGITOS (11 DOWNTO 8);
							DIGITOS (11 DOWNTO 8) = DIGITOS (7 DOWNTO 4);
							DIGITOS (7 DOWNTO 4) = DIGITOS (3 DOWNTO 0);
							DIGITOS (3 DOWNTO 0) = ENTRADA;
							COUNT := COUNT + 1
					END CASE;
				END IF;
		END CASE;

	END PROCESS;

	RESETN <= KEY(0);

	pwn: PWN PORT MAP (
		CLOCK, RESET, ENABLE, DUTY,
		COUT
	);

	dig_calc: conv_calc PORT MAP (
		key0(7 DOWNTO 0), ENTRADA
	);

	somador0: somadorBinarioParalelo PORT MAP (
		A (3 DOWNTO 0), B (3 DOWNTO 0), 0,
		DBUFFER (3 DOWNTO 0), C(0)
	);
	somador1: somadorBinarioParalelo PORT MAP (
		A (7 DOWNTO 4), B (7 DOWNTO 4), C(0),
		DBUFFER (7 DOWNTO 4), C(1)
	);
	somador2: somadorBinarioParalelo PORT MAP (
		A (11 DOWNTO 8), B (11 DOWNTO 8), C(1),
		DBUFFER (7 DOWNTO 4), C(2)
	);
	somador3: somadorBinarioParalelo PORT MAP (
		A (15 DOWNTO 12), B (15 DOWNTO 12), C(2),
		DBUFFER (7 DOWNTO 4), C(3)
	);

	hexseg0: conv_7seg PORT MAP (
		DIGITOS (3 DOWNTO 0), HEX0
	);
	hexseg1: conv_7seg PORT MAP (
		DIGITOS (7 DOWNTO 4), HEX1
	);
	hexseg2: conv_7seg PORT MAP (
		DIGITOS (11 DOWNTO 8), HEX2
	);
	hexseg3: conv_7seg PORT MAP (
		DIGITOS (15 DOWNTO 12), HEX3
	);

	kbd_ctrl : kbdex_ctrl GENERIC MAP(24000) PORT MAP(
		PS2_DAT, PS2_CLK, CLOCK_24(0), KEY(1), resetn, lights(1) & lights(2) & lights(0),
		key_on, key_code(15 DOWNTO 0) => key0
	);

END funcionamento;